`timescale 1ps/1ps

module mux_16to1_tb;
    reg [15:0] t_datain;
	reg [3:0] t_select;
	wire t_outd;
    
    mux_16to1 dut1 (.datain(t_datain), .select(t_select), .outd(t_outd));

    initial begin
        #0 
        t_datain = 0; 
        t_select = 0;
    end

    initial begin
        // 0
        #10 t_datain = 1;
        #10 t_select = 0;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 1
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 2
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 3
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 4
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 5
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 6
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 7
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 8
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 9
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 10
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 11
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 12
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 13
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 14
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // 15
        t_datain = t_datain << 1;
        #10 t_select = 1;
        #10 t_select = 2;
        #10 t_select = 3;
        #10 t_select = 4;
        #10 t_select = 5;
        #10 t_select = 6;
        #10 t_select = 7;
        #10 t_select = 8;
        #10 t_select = 9;
        #10 t_select = 10;
        #10 t_select = 11;
        #10 t_select = 12;
        #10 t_select = 13;
        #10 t_select = 14;
        #10 t_select = 15;
        #10 t_select = 0;
        // spacial
        #10 t_select = 4'b000x;
        #10 t_select = 4'b00xx;
        #10 t_select = 4'b000z;
        #10 t_select = 4'b00zz;
        #10 t_select = 4'b00xz;
        #10 t_select = 4'b00zx;
        #10 t_select = 4'bxxxx;
        $stop;
    end
endmodule